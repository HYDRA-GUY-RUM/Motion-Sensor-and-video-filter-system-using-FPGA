module Color_Detector_FSM(clk,	data,	startofpacket,	endofpacket, right, up, left, down, LEDR);

	input clk, startofpacket,	endofpacket;
	input [29:0]data;
	output right, up, left, down;
	output [7:0]LEDR;
	reg a, b, c, d, z, k, a1, b1, c1, d1, z1, k1;

		always @(*)						
		begin		
		//This is where all the cases are executed 
			if(startofpacket == 1)
			begin
			//This is executed only when we want to start reading a frame 
				z1=0;
				a1=0;
				b1=0;
				c1=0;
				d1=0;
				k1=1;
			end
			if(endofpacket == 1)
			begin
			//This is executed when we have finished reading a frame 
				k1=0;
			end
		end
			
		always @(posedge clk)	
		begin
		a = a1;
		b = b1;
		c = c1;
		d = d1;
		z = z1;
		k = k1;
			if(k==1)
			begin
			//We read data when k = 1
					if(data[9:0] > 10'b1001011000 && data[19:10] > 10'b1001011000 && data[29:20] > 10'b1001011000)
					begin
					//This is executed only when the color of the pixel is white(ie. above R[600], G[600] and B[600])
						if((z >= 320 && z < 640)
							 || (z >= 960 && z < 1280)
							 || (z >= 1600 && z < 1920)
							 || (z >= 2240 && z < 2560)
							 || (z >= 2880 && z < 3200)
							 || (z >= 3520 && z < 3840)
							 || (z >= 4160 && z < 4480)
							 || (z >= 4800 && z < 5120)
							 || (z >= 5440 && z < 5760)
							 || (z >= 6080 && z < 6400)
							 || (z >= 6720 && z < 7040)
							 || (z >= 7360 && z < 7680)
							 || (z >= 8000 && z < 8320)
							 || (z >= 8640 && z < 8960)
							 || (z >= 9280 && z < 9600)
							 || (z >= 9920 && z < 10240)
							 || (z >= 10560 && z < 10880)
							 || (z >= 11200 && z < 11520)
							 || (z >= 11840 && z < 12160)
							 || (z >= 12480 && z < 12800)
							 || (z >= 13120 && z < 13440)
							 || (z >= 13760 && z < 14080)
							 || (z >= 14400 && z < 14720)
							 || (z >= 15040 && z < 15360)
							 || (z >= 15680 && z < 16000)
							 || (z >= 16320 && z < 16640)
							 || (z >= 16960 && z < 17280)
							 || (z >= 17600 && z < 17920)
							 || (z >= 18240 && z < 18560)
							 || (z >= 18880 && z < 19200)
							 || (z >= 19520 && z < 19840)
							 || (z >= 20160 && z < 20480)
							 || (z >= 20800 && z < 21120)
							 || (z >= 21440 && z < 21760)
							 || (z >= 22080 && z < 22400)
							 || (z >= 22720 && z < 23040)
							 || (z >= 23360 && z < 23680)
							 || (z >= 24000 && z < 24320)
							 || (z >= 24640 && z < 24960)
							 || (z >= 25280 && z < 25600)
							 || (z >= 25920 && z < 26240)
							 || (z >= 26560 && z < 26880)
							 || (z >= 27200 && z < 27520)
							 || (z >= 27840 && z < 28160)
							 || (z >= 28480 && z < 28800)
							 || (z >= 29120 && z < 29440)
							 || (z >= 29760 && z < 30080)
							 || (z >= 30400 && z < 30720)
							 || (z >= 31040 && z < 31360)
							 || (z >= 31680 && z < 32000)
							 || (z >= 32320 && z < 32640)
							 || (z >= 32960 && z < 33280)
							 || (z >= 33600 && z < 33920)
							 || (z >= 34240 && z < 34560)
							 || (z >= 34880 && z < 35200)
							 || (z >= 35520 && z < 35840)
							 || (z >= 36160 && z < 36480)
							 || (z >= 36800 && z < 37120)
							 || (z >= 37440 && z < 37760)
							 || (z >= 38080 && z < 38400)
							 || (z >= 38720 && z < 39040)
							 || (z >= 39360 && z < 39680)
							 || (z >= 40000 && z < 40320)
							 || (z >= 40640 && z < 40960)
							 || (z >= 41280 && z < 41600)
							 || (z >= 41920 && z < 42240)
							 || (z >= 42560 && z < 42880)
							 || (z >= 43200 && z < 43520)
							 || (z >= 43840 && z < 44160)
							 || (z >= 44480 && z < 44800)
							 || (z >= 45120 && z < 45440)
							 || (z >= 45760 && z < 46080)
							 || (z >= 46400 && z < 46720)
							 || (z >= 47040 && z < 47360)
							 || (z >= 47680 && z < 48000)
							 || (z >= 48320 && z < 48640)
							 || (z >= 48960 && z < 49280)
							 || (z >= 49600 && z < 49920)
							 || (z >= 50240 && z < 50560)
							 || (z >= 50880 && z < 51200)
							 || (z >= 51520 && z < 51840)
							 || (z >= 52160 && z < 52480)
							 || (z >= 52800 && z < 53120)
							 || (z >= 53440 && z < 53760)
							 || (z >= 54080 && z < 54400)
							 || (z >= 54720 && z < 55040)
							 || (z >= 55360 && z < 55680)
							 || (z >= 56000 && z < 56320)
							 || (z >= 56640 && z < 56960)
							 || (z >= 57280 && z < 57600)
							 || (z >= 57920 && z < 58240)
							 || (z >= 58560 && z < 58880)
							 || (z >= 59200 && z < 59520)
							 || (z >= 59840 && z < 60160)
							 || (z >= 60480 && z < 60800)
							 || (z >= 61120 && z < 61440)
							 || (z >= 61760 && z < 62080)
							 || (z >= 62400 && z < 62720)
							 || (z >= 63040 && z < 63360)
							 || (z >= 63680 && z < 64000)
							 || (z >= 64320 && z < 64640)
							 || (z >= 64960 && z < 65280)
							 || (z >= 65600 && z < 65920)
							 || (z >= 66240 && z < 66560)
							 || (z >= 66880 && z < 67200)
							 || (z >= 67520 && z < 67840)
							 || (z >= 68160 && z < 68480)
							 || (z >= 68800 && z < 69120)
							 || (z >= 69440 && z < 69760)
							 || (z >= 70080 && z < 70400)
							 || (z >= 70720 && z < 71040)
							 || (z >= 71360 && z < 71680)
							 || (z >= 72000 && z < 72320)
							 || (z >= 72640 && z < 72960)
							 || (z >= 73280 && z < 73600)
							 || (z >= 73920 && z < 74240)
							 || (z >= 74560 && z < 74880)
							 || (z >= 75200 && z < 75520)
							 || (z >= 75840 && z < 76160)
							 || (z >= 76480 && z < 76800)
							 || (z >= 77120 && z < 77440)
							 || (z >= 77760 && z < 78080)
							 || (z >= 78400 && z < 78720)
							 || (z >= 79040 && z < 79360)
							 || (z >= 79680 && z < 80000)
							 || (z >= 80320 && z < 80640)
							 || (z >= 80960 && z < 81280)
							 || (z >= 81600 && z < 81920)
							 || (z >= 82240 && z < 82560)
							 || (z >= 82880 && z < 83200)
							 || (z >= 83520 && z < 83840)
							 || (z >= 84160 && z < 84480)
							 || (z >= 84800 && z < 85120)
							 || (z >= 85440 && z < 85760)
							 || (z >= 86080 && z < 86400)
							 || (z >= 86720 && z < 87040)
							 || (z >= 87360 && z < 87680)
							 || (z >= 88000 && z < 88320)
							 || (z >= 88640 && z < 88960)
							 || (z >= 89280 && z < 89600)
							 || (z >= 89920 && z < 90240)
							 || (z >= 90560 && z < 90880)
							 || (z >= 91200 && z < 91520)
							 || (z >= 91840 && z < 92160)
							 || (z >= 92480 && z < 92800)
							 || (z >= 93120 && z < 93440)
							 || (z >= 93760 && z < 94080)
							 || (z >= 94400 && z < 94720)
							 || (z >= 95040 && z < 95360)
							 || (z >= 95680 && z < 96000)
							 || (z >= 96320 && z < 96640)
							 || (z >= 96960 && z < 97280)
							 || (z >= 97600 && z < 97920)
							 || (z >= 98240 && z < 98560)
							 || (z >= 98880 && z < 99200)
							 || (z >= 99520 && z < 99840)
							 || (z >= 100160 && z < 100480)
							 || (z >= 100800 && z < 101120)
							 || (z >= 101440 && z < 101760)
							 || (z >= 102080 && z < 102400)
							 || (z >= 102720 && z < 103040)
							 || (z >= 103360 && z < 103680)
							 || (z >= 104000 && z < 104320)
							 || (z >= 104640 && z < 104960)
							 || (z >= 105980 && z < 105600)
							 || (z >= 105920 && z < 106240)
							 || (z >= 106560 && z < 106880)
							 || (z >= 107200 && z < 107520)
							 || (z >= 107840 && z < 108160)
							 || (z >= 108480 && z < 108800)
							 || (z >= 109120 && z < 109440)
							 || (z >= 109760 && z < 110080)
							 || (z >= 110400 && z < 110720)
							 || (z >= 111040 && z < 111360)
							 || (z >= 111680 && z < 112000)
							 || (z >= 112320 && z < 112640)
							 || (z >= 112960 && z < 113280)
							 || (z >= 113600 && z < 113920)
							 || (z >= 114240 && z < 114560)
							 || (z >= 114880 && z < 115200)
							 || (z >= 115520 && z < 115840)
							 || (z >= 116160 && z < 116480)
							 || (z >= 116800 && z < 117120)
							 || (z >= 117440 && z < 117760)
							 || (z >= 118080 && z < 118400)
							 || (z >= 118720 && z < 119040)
							 || (z >= 119360 && z < 119680)
							 || (z >= 120000 && z < 120320)
							 || (z >= 120640 && z < 120960)
							 || (z >= 121280 && z < 121600)
							 || (z >= 121920 && z < 122240)
							 || (z >= 122560 && z < 122880)
							 || (z >= 123200 && z < 123520)
							 || (z >= 123840 && z < 124160)
							 || (z >= 124480 && z < 124800)
							 || (z >= 125120 && z < 125440)
							 || (z >= 125760 && z < 126080)
							 || (z >= 126040 && z < 126720)
							 || (z >= 127040 && z < 127360)
							 || (z >= 127680 && z < 128000)
							 || (z >= 128320 && z < 128640)
							 || (z >= 128960 && z < 129280)
							 || (z >= 129600 && z < 129920)
							 || (z >= 130240 && z < 130560)
							 || (z >= 130880 && z < 131200)
							 || (z >= 131520 && z < 131840)
							 || (z >= 132160 && z < 132480)
							 || (z >= 132800 && z < 133120)
							 || (z >= 133440 && z < 133760)
							 || (z >= 134080 && z < 134400)
							 || (z >= 134720 && z < 135040)
							 || (z >= 135360 && z < 135680)
							 || (z >= 136000 && z < 136320)
							 || (z >= 136640 && z < 136960)
							 || (z >= 137280 && z < 137600)
							 || (z >= 137920 && z < 138240)
							 || (z >= 138560 && z < 138880)
							 || (z >= 139200 && z < 139520)
							 || (z >= 139840 && z < 140160)
							 || (z >= 140480 && z < 140800)
							 || (z >= 141121 && z < 141440)
							 || (z >= 141760 && z < 142080)
							 || (z >= 142400 && z < 142720)
							 || (z >= 143040 && z < 143360)
							 || (z >= 143680 && z < 144000)
							 || (z >= 144320 && z < 144640)
							 || (z >= 144960 && z < 145280)
							 || (z >= 145600 && z < 145920)
							 || (z >= 146240 && z < 146560)
							 || (z >= 146880 && z < 147200)
							 || (z >= 147520 && z < 147840)
							 || (z >= 148160 && z < 148480)
							 || (z >= 148800 && z < 149120)
							 || (z >= 149440 && z < 149760)
							 || (z >= 150080 && z < 150400)
							 || (z >= 150720 && z < 151040)
							 || (z >= 151360 && z < 151680)
							 || (z >= 152000 && z < 152320)
							 || (z >= 152640 && z < 152960)
							 || (z >= 153280 && z < 153600)
							 || (z >= 153920 && z < 154240)
							 || (z >= 154560 && z < 154880)
							 || (z >= 155200 && z < 155520)
							 || (z >= 155840 && z < 156160)
							 || (z >= 156480 && z < 156800)
							 || (z >= 157120 && z < 157440)
							 || (z >= 157760 && z < 158080)
							 || (z >= 158400 && z < 158720)
							 || (z >= 159040 && z < 159360)
							 || (z >= 159680 && z < 160000)
							 || (z >= 160320 && z < 160640)
							 || (z >= 160960 && z < 161280)
							 || (z >= 161600 && z < 161920)
							 || (z >= 162240 && z < 162560)
							 || (z >= 162880 && z < 163200)
							 || (z >= 163520 && z < 163840)
							 || (z >= 164160 && z < 164480)
							 || (z >= 164800 && z < 165120)
							 || (z >= 165440 && z < 165760)
							 || (z >= 166080 && z < 166400)
							 || (z >= 166720 && z < 167040)
							 || (z >= 167360 && z < 167680)
							 || (z >= 168000 && z < 168320)
							 || (z >= 168640 && z < 168960)
							 || (z >= 169280 && z < 169600)
							 || (z >= 169920 && z < 170240)
							 || (z >= 170560 && z < 170880)
							 || (z >= 171200 && z < 171520)
							 || (z >= 171840 && z < 172160)
							 || (z >= 172480 && z < 172800)
							 || (z >= 173120 && z < 173440)
							 || (z >= 173760 && z < 174080)
							 || (z >= 174400 && z < 174720)
							 || (z >= 175040 && z < 175360)
							 || (z >= 175680 && z < 176000)
							 || (z >= 176320 && z < 176640)
							 || (z >= 176960 && z < 177280)
							 || (z >= 177600 && z < 177920)
							 || (z >= 178240 && z < 178560)
							 || (z >= 178880 && z < 179200)
							 || (z >= 179520 && z < 179840)
							 || (z >= 180160 && z < 180480)
							 || (z >= 180800 && z < 181120)
							 || (z >= 181440 && z < 181760)
							 || (z >= 182080 && z < 182400)
							 || (z >= 182720 && z < 183040)
							 || (z >= 183360 && z < 183680)
							 || (z >= 184000 && z < 184320)
							 || (z >= 184640 && z < 184960)
							 || (z >= 185280 && z < 185600)
							 || (z >= 185920 && z < 186240)
							 || (z >= 186560 && z < 186880)
							 || (z >= 187200 && z < 187520)
							 || (z >= 187840 && z < 188160)
							 || (z >= 188480 && z < 188800)
							 || (z >= 189120 && z < 189440)
							 || (z >= 189760 && z < 190080)
							 || (z >= 190400 && z < 190720)
							 || (z >= 191040 && z < 191360)
							 || (z >= 191680 && z < 192000)
							 || (z >= 192320 && z < 192640)
							 || (z >= 192960 && z < 193280)
							 || (z >= 193600 && z < 193920)
							 || (z >= 194240 && z < 194560)
							 || (z >= 194880 && z < 195200)
							 || (z >= 195520 && z < 195840)
							 || (z >= 196160 && z < 196480)
							 || (z >= 196800 && z < 197120)
							 || (z >= 197440 && z < 197760)
							 || (z >= 198080 && z < 198400)
							 || (z >= 198720 && z < 199040)
							 || (z >= 199360 && z < 199680)
							 || (z >= 200000 && z < 200320)
							 || (z >= 200640 && z < 200960)
							 || (z >= 201280 && z < 201600)
							 || (z >= 201920 && z < 202240)
							 || (z >= 202560 && z < 202880)
							 || (z >= 203200 && z < 203520)
							 || (z >= 203840 && z < 204160)
							 || (z >= 204480 && z < 204800)
							 || (z >= 205120 && z < 205440)
							 || (z >= 205760 && z < 206080)
							 || (z >= 206400 && z < 206720)
							 || (z >= 207040 && z < 207360)
							 || (z >= 207680 && z < 208000)
							 || (z >= 208320 && z < 208640)
							 || (z >= 208960 && z < 209280)
							 || (z >= 209600 && z < 209320)
							 || (z >= 210240 && z < 210560)
							 || (z >= 210880 && z < 211200)
							 || (z >= 211520 && z < 211840)
							 || (z >= 212160 && z < 212480)
							 || (z >= 212800 && z < 213120)
							 || (z >= 213440 && z < 213760)
							 || (z >= 214080 && z < 214400)
							 || (z >= 214720 && z < 215040)
							 || (z >= 215360 && z < 215680)
							 || (z >= 216000 && z < 216320)
							 || (z >= 216640 && z < 216960)
							 || (z >= 217280 && z < 217600)
							 || (z >= 217920 && z < 218240)
							 || (z >= 218560 && z < 218880)
							 || (z >= 219200 && z < 219520)
							 || (z >= 219840 && z < 220160)
							 || (z >= 220480 && z < 220800)
							 || (z >= 221120 && z < 221440)
							 || (z >= 221760 && z < 222080)
							 || (z >= 222400 && z < 222720)
							 || (z >= 223040 && z < 223360)
							 || (z >= 223680 && z < 224000)
							 || (z >= 224320 && z < 224640)
							 || (z >= 224960 && z < 225280)
							 || (z >= 225600 && z < 225920)
							 || (z >= 226240 && z < 226560)
							 || (z >= 226880 && z < 227200)
							 || (z >= 227520 && z < 227840)
							 || (z >= 228160 && z < 228480)
							 || (z >= 228800 && z < 229120)
							 || (z >= 229440 && z < 229760)
							 || (z >= 230080 && z < 230400)
							 || (z >= 230720 && z < 231040)
							 || (z >= 231360 && z < 231680)
							 || (z >= 232000 && z < 232320)
							 || (z >= 232640 && z < 232960)
							 || (z >= 233280 && z < 233600)
							 || (z >= 233920 && z < 234240)
							 || (z >= 234560 && z < 234880)
							 || (z >= 235200 && z < 235520)
							 || (z >= 235840 && z < 236160)
							 || (z >= 236480 && z < 236800)
							 || (z >= 237120 && z < 237440)
							 || (z >= 237760 && z < 238080)
							 || (z >= 238400 && z < 238720)
							 || (z >= 239040 && z < 239360)
							 || (z >= 239680 && z < 240000)
							 || (z >= 240320 && z < 240640)
							 || (z >= 240960 && z < 241280)
							 || (z >= 241600 && z < 241920)
							 || (z >= 242240 && z < 242560)
							 || (z >= 242880 && z < 243200)
							 || (z >= 243520 && z < 243840)
							 || (z >= 244160 && z < 244480)
							 || (z >= 244800 && z < 245120)
							 || (z >= 245440 && z < 245760)
							 || (z >= 246080 && z < 246400)
							 || (z >= 246720 && z < 247040)
							 || (z >= 247360 && z < 247680)
							 || (z >= 248000 && z < 248320)
							 || (z >= 248640 && z < 248960)
							 || (z >= 249280 && z < 249600)
							 || (z >= 249920 && z < 250240)
							 || (z >= 250560 && z < 250880)
							 || (z >= 251200 && z < 251520)
							 || (z >= 251840 && z < 252160)
							 || (z >= 252480 && z < 252800)
							 || (z >= 253120 && z < 253440)
							 || (z >= 253760 && z < 254080)
							 || (z >= 254400 && z < 254720)
							 || (z >= 255040 && z < 255360)
							 || (z >= 255680 && z < 256000)
							 || (z >= 256320 && z < 256640)
							 || (z >= 256960 && z < 257280)
							 || (z >= 257600 && z < 257920)
							 || (z >= 258240 && z < 258560)
							 || (z >= 258880 && z < 259200)
							 || (z >= 259520 && z < 259840)
							 || (z >= 260160 && z < 260480)
							 || (z >= 260800 && z < 261120)
							 || (z >= 261440 && z < 261760)
							 || (z >= 262080 && z < 262400)
							 || (z >= 262720 && z < 263040)
							 || (z >= 263360 && z < 236680)
							 || (z >= 264000 && z < 264320)
							 || (z >= 264640 && z < 264960)
							 || (z >= 265280 && z < 265600)
							 || (z >= 265920 && z < 266240)
							 || (z >= 266560 && z < 266880)
							 || (z >= 267200 && z < 267520)
							 || (z >= 267840 && z < 268160)
							 || (z >= 268480 && z < 268800)
							 || (z >= 269120 && z < 269440)
							 || (z >= 269760 && z < 270080)
							 || (z >= 270400 && z < 270720)
							 || (z >= 271040 && z < 271360)
							 || (z >= 271680 && z < 272000)
							 || (z >= 272320 && z < 272640)
							 || (z >= 272960 && z < 273280)
							 || (z >= 273600 && z < 273920)
							 || (z >= 272240 && z < 274560)
							 || (z >= 274880 && z < 275200)
							 || (z >= 275520 && z < 275840)
							 || (z >= 276160 && z < 276480)
							 || (z >= 276800 && z < 277120)
							 || (z >= 277440 && z < 277760)
							 || (z >= 278080 && z < 278400)
							 || (z >= 278720 && z < 279040)
							 || (z >= 279360 && z < 279680)
							 || (z >= 280000 && z < 280320)
							 || (z >= 280640 && z < 280960)
							 || (z >= 281280 && z < 281600)
							 || (z >= 281920 && z < 282240)
							 || (z >= 282560 && z < 282880)
							 || (z >= 283200 && z < 283520)
							 || (z >= 283840 && z < 284160)
							 || (z >= 284480 && z < 284800)
							 || (z >= 285120 && z < 285440)
							 || (z >= 285760 && z < 286080)
							 || (z >= 286400 && z < 286720)
							 || (z >= 287040 && z < 287360)
							 || (z >= 287680 && z < 288000)
							 || (z >= 288320 && z < 288640)
							 || (z >= 288960 && z < 289280)
							 || (z >= 289600 && z < 289920)
							 || (z >= 290240 && z < 290560)
							 || (z >= 290880 && z < 291200)
							 || (z >= 291520 && z < 291840)
							 || (z >= 292160 && z < 292480)
							 || (z >= 292800 && z < 293120)
							 || (z >= 293440 && z < 293760)
							 || (z >= 294080 && z < 294400)
							 || (z >= 294720 && z < 295040)
							 || (z >= 295360 && z < 295680)
							 || (z >= 296000 && z < 296320)
							 || (z >= 296640 && z < 296960)
							 || (z >= 297280 && z < 297600)
							 || (z >= 297920 && z < 298240)
							 || (z >= 298560 && z < 298880)
							 || (z >= 299200 && z < 299520)
							 || (z >= 299840 && z < 300160)
							 || (z >= 300480 && z < 300800)
							 || (z >= 301120 && z < 301440)
							 || (z >= 301760 && z < 302080)
							 || (z >= 302400 && z < 302720)
							 || (z >= 303040 && z < 303360)
							 || (z >= 303680 && z < 304000)
							 || (z >= 304320 && z < 304640)
							 || (z >= 304960 && z < 305280)
							 || (z >= 305600 && z < 305920)
							 || (z >= 306240 && z < 306560)
							 || (z >= 306880 && z < 307200))
						begin
						//This is executed when the white pixel belongs to the right half(a direction)
							a=a+1;
						end
						if(z >= 0 && z < 153600)
						begin
						//This is executed when the white pixel belongs to the upper half(b direction)
							b = b+1;
						end
						if((z >= (-320) + 320 && z < (-320) + 640)
							 || (z >= (-320) + 960 && z < (-320) + 1280)
							 || (z >= (-320) + 1600 && z < (-320) + 1920)
							 || (z >= (-320) + 2240 && z < (-320) + 2560)
							 || (z >= (-320) + 2880 && z < (-320) + 3200)
							 || (z >= (-320) + 3520 && z < (-320) + 3840)
							 || (z >= (-320) + 4160 && z < (-320) + 4480)
							 || (z >= (-320) + 4800 && z < (-320) + 5120)
							 || (z >= (-320) + 5440 && z < (-320) + 5760)
							 || (z >= (-320) + 6080 && z < (-320) + 6400)
							 || (z >= (-320) + 6720 && z < (-320) + 7040)
							 || (z >= (-320) + 7360 && z < (-320) + 7680)
							 || (z >= (-320) + 8000 && z < (-320) + 8320)
							 || (z >= (-320) + 8640 && z < (-320) + 8960)
							 || (z >= (-320) + 9280 && z < (-320) + 9600)
							 || (z >= (-320) + 9920 && z < (-320) + 10240)
							 || (z >= (-320) + 10560 && z < (-320) + 10880)
							 || (z >= (-320) + 11200 && z < (-320) + 11520)
							 || (z >= (-320) + 11840 && z < (-320) + 12160)
							 || (z >= (-320) + 12480 && z < (-320) + 12800)
							 || (z >= (-320) + 13120 && z < (-320) + 13440)
							 || (z >= (-320) + 13760 && z < (-320) + 14080)
							 || (z >= (-320) + 14400 && z < (-320) + 14720)
							 || (z >= (-320) + 15040 && z < (-320) + 15360)
							 || (z >= (-320) + 15680 && z < (-320) + 16000)
							 || (z >= (-320) + 16320 && z < (-320) + 16640)
							 || (z >= (-320) + 16960 && z < (-320) + 17280)
							 || (z >= (-320) + 17600 && z < (-320) + 17920)
							 || (z >= (-320) + 18240 && z < (-320) + 18560)
							 || (z >= (-320) + 18880 && z < (-320) + 19200)
							 || (z >= (-320) + 19520 && z < (-320) + 19840)
							 || (z >= (-320) + 20160 && z < (-320) + 20480)
							 || (z >= (-320) + 20800 && z < (-320) + 21120)
							 || (z >= (-320) + 21440 && z < (-320) + 21760)
							 || (z >= (-320) + 22080 && z < (-320) + 22400)
							 || (z >= (-320) + 22720 && z < (-320) + 23040)
							 || (z >= (-320) + 23360 && z < (-320) + 23680)
							 || (z >= (-320) + 24000 && z < (-320) + 24320)
							 || (z >= (-320) + 24640 && z < (-320) + 24960)
							 || (z >= (-320) + 25280 && z < (-320) + 25600)
							 || (z >= (-320) + 25920 && z < (-320) + 26240)
							 || (z >= (-320) + 26560 && z < (-320) + 26880)
							 || (z >= (-320) + 27200 && z < (-320) + 27520)
							 || (z >= (-320) + 27840 && z < (-320) + 28160)
							 || (z >= (-320) + 28480 && z < (-320) + 28800)
							 || (z >= (-320) + 29120 && z < (-320) + 29440)
							 || (z >= (-320) + 29760 && z < (-320) + 30080)
							 || (z >= (-320) + 30400 && z < (-320) + 30720)
							 || (z >= (-320) + 31040 && z < (-320) + 31360)
							 || (z >= (-320) + 31680 && z < (-320) + 32000)
							 || (z >= (-320) + 32320 && z < (-320) + 32640)
							 || (z >= (-320) + 32960 && z < (-320) + 33280)
							 || (z >= (-320) + 33600 && z < (-320) + 33920)
							 || (z >= (-320) + 34240 && z < (-320) + 34560)
							 || (z >= (-320) + 34880 && z < (-320) + 35200)
							 || (z >= (-320) + 35520 && z < (-320) + 35840)
							 || (z >= (-320) + 36160 && z < (-320) + 36480)
							 || (z >= (-320) + 36800 && z < (-320) + 37120)
							 || (z >= (-320) + 37440 && z < (-320) + 37760)
							 || (z >= (-320) + 38080 && z < (-320) + 38400)
							 || (z >= (-320) + 38720 && z < (-320) + 39040)
							 || (z >= (-320) + 39360 && z < (-320) + 39680)
							 || (z >= (-320) + 40000 && z < (-320) + 40320)
							 || (z >= (-320) + 40640 && z < (-320) + 40960)
							 || (z >= (-320) + 41280 && z < (-320) + 41600)
							 || (z >= (-320) + 41920 && z < (-320) + 42240)
							 || (z >= (-320) + 42560 && z < (-320) + 42880)
							 || (z >= (-320) + 43200 && z < (-320) + 43520)
							 || (z >= (-320) + 43840 && z < (-320) + 44160)
							 || (z >= (-320) + 44480 && z < (-320) + 44800)
							 || (z >= (-320) + 45120 && z < (-320) + 45440)
							 || (z >= (-320) + 45760 && z < (-320) + 46080)
							 || (z >= (-320) + 46400 && z < (-320) + 46720)
							 || (z >= (-320) + 47040 && z < (-320) + 47360)
							 || (z >= (-320) + 47680 && z < (-320) + 48000)
							 || (z >= (-320) + 48320 && z < (-320) + 48640)
							 || (z >= (-320) + 48960 && z < (-320) + 49280)
							 || (z >= (-320) + 49600 && z < (-320) + 49920)
							 || (z >= (-320) + 50240 && z < (-320) + 50560)
							 || (z >= (-320) + 50880 && z < (-320) + 51200)
							 || (z >= (-320) + 51520 && z < (-320) + 51840)
							 || (z >= (-320) + 52160 && z < (-320) + 52480)
							 || (z >= (-320) + 52800 && z < (-320) + 53120)
							 || (z >= (-320) + 53440 && z < (-320) + 53760)
							 || (z >= (-320) + 54080 && z < (-320) + 54400)
							 || (z >= (-320) + 54720 && z < (-320) + 55040)
							 || (z >= (-320) + 55360 && z < (-320) + 55680)
							 || (z >= (-320) + 56000 && z < (-320) + 56320)
							 || (z >= (-320) + 56640 && z < (-320) + 56960)
							 || (z >= (-320) + 57280 && z < (-320) + 57600)
							 || (z >= (-320) + 57920 && z < (-320) + 58240)
							 || (z >= (-320) + 58560 && z < (-320) + 58880)
							 || (z >= (-320) + 59200 && z < (-320) + 59520)
							 || (z >= (-320) + 59840 && z < (-320) + 60160)
							 || (z >= (-320) + 60480 && z < (-320) + 60800)
							 || (z >= (-320) + 61120 && z < (-320) + 61440)
							 || (z >= (-320) + 61760 && z < (-320) + 62080)
							 || (z >= (-320) + 62400 && z < (-320) + 62720)
							 || (z >= (-320) + 63040 && z < (-320) + 63360)
							 || (z >= (-320) + 63680 && z < (-320) + 64000)
							 || (z >= (-320) + 64320 && z < (-320) + 64640)
							 || (z >= (-320) + 64960 && z < (-320) + 65280)
							 || (z >= (-320) + 65600 && z < (-320) + 65920)
							 || (z >= (-320) + 66240 && z < (-320) + 66560)
							 || (z >= (-320) + 66880 && z < (-320) + 67200)
							 || (z >= (-320) + 67520 && z < (-320) + 67840)
							 || (z >= (-320) + 68160 && z < (-320) + 68480)
							 || (z >= (-320) + 68800 && z < (-320) + 69120)
							 || (z >= (-320) + 69440 && z < (-320) + 69760)
							 || (z >= (-320) + 70080 && z < (-320) + 70400)
							 || (z >= (-320) + 70720 && z < (-320) + 71040)
							 || (z >= (-320) + 71360 && z < (-320) + 71680)
							 || (z >= (-320) + 72000 && z < (-320) + 72320)
							 || (z >= (-320) + 72640 && z < (-320) + 72960)
							 || (z >= (-320) + 73280 && z < (-320) + 73600)
							 || (z >= (-320) + 73920 && z < (-320) + 74240)
							 || (z >= (-320) + 74560 && z < (-320) + 74880)
							 || (z >= (-320) + 75200 && z < (-320) + 75520)
							 || (z >= (-320) + 75840 && z < (-320) + 76160)
							 || (z >= (-320) + 76480 && z < (-320) + 76800)
							 || (z >= (-320) + 77120 && z < (-320) + 77440)
							 || (z >= (-320) + 77760 && z < (-320) + 78080)
							 || (z >= (-320) + 78400 && z < (-320) + 78720)
							 || (z >= (-320) + 79040 && z < (-320) + 79360)
							 || (z >= (-320) + 79680 && z < (-320) + 80000)
							 || (z >= (-320) + 80320 && z < (-320) + 80640)
							 || (z >= (-320) + 80960 && z < (-320) + 81280)
							 || (z >= (-320) + 81600 && z < (-320) + 81920)
							 || (z >= (-320) + 82240 && z < (-320) + 82560)
							 || (z >= (-320) + 82880 && z < (-320) + 83200)
							 || (z >= (-320) + 83520 && z < (-320) + 83840)
							 || (z >= (-320) + 84160 && z < (-320) + 84480)
							 || (z >= (-320) + 84800 && z < (-320) + 85120)
							 || (z >= (-320) + 85440 && z < (-320) + 85760)
							 || (z >= (-320) + 86080 && z < (-320) + 86400)
							 || (z >= (-320) + 86720 && z < (-320) + 87040)
							 || (z >= (-320) + 87360 && z < (-320) + 87680)
							 || (z >= (-320) + 88000 && z < (-320) + 88320)
							 || (z >= (-320) + 88640 && z < (-320) + 88960)
							 || (z >= (-320) + 89280 && z < (-320) + 89600)
							 || (z >= (-320) + 89920 && z < (-320) + 90240)
							 || (z >= (-320) + 90560 && z < (-320) + 90880)
							 || (z >= (-320) + 91200 && z < (-320) + 91520)
							 || (z >= (-320) + 91840 && z < (-320) + 92160)
							 || (z >= (-320) + 92480 && z < (-320) + 92800)
							 || (z >= (-320) + 93120 && z < (-320) + 93440)
							 || (z >= (-320) + 93760 && z < (-320) + 94080)
							 || (z >= (-320) + 94400 && z < (-320) + 94720)
							 || (z >= (-320) + 95040 && z < (-320) + 95360)
							 || (z >= (-320) + 95680 && z < (-320) + 96000)
							 || (z >= (-320) + 96320 && z < (-320) + 96640)
							 || (z >= (-320) + 96960 && z < (-320) + 97280)
							 || (z >= (-320) + 97600 && z < (-320) + 97920)
							 || (z >= (-320) + 98240 && z < (-320) + 98560)
							 || (z >= (-320) + 98880 && z < (-320) + 99200)
							 || (z >= (-320) + 99520 && z < (-320) + 99840)
							 || (z >= (-320) + 100160 && z < (-320) + 100480)
							 || (z >= (-320) + 100800 && z < (-320) + 101120)
							 || (z >= (-320) + 101440 && z < (-320) + 101760)
							 || (z >= (-320) + 102080 && z < (-320) + 102400)
							 || (z >= (-320) + 102720 && z < (-320) + 103040)
							 || (z >= (-320) + 103360 && z < (-320) + 103680)
							 || (z >= (-320) + 104000 && z < (-320) + 104320)
							 || (z >= (-320) + 104640 && z < (-320) + 104960)
							 || (z >= (-320) + 105980 && z < (-320) + 105600)
							 || (z >= (-320) + 105920 && z < (-320) + 106240)
							 || (z >= (-320) + 106560 && z < (-320) + 106880)
							 || (z >= (-320) + 107200 && z < (-320) + 107520)
							 || (z >= (-320) + 107840 && z < (-320) + 108160)
							 || (z >= (-320) + 108480 && z < (-320) + 108800)
							 || (z >= (-320) + 109120 && z < (-320) + 109440)
							 || (z >= (-320) + 109760 && z < (-320) + 110080)
							 || (z >= (-320) + 110400 && z < (-320) + 110720)
							 || (z >= (-320) + 111040 && z < (-320) + 111360)
							 || (z >= (-320) + 111680 && z < (-320) + 112000)
							 || (z >= (-320) + 112320 && z < (-320) + 112640)
							 || (z >= (-320) + 112960 && z < (-320) + 113280)
							 || (z >= (-320) + 113600 && z < (-320) + 113920)
							 || (z >= (-320) + 114240 && z < (-320) + 114560)
							 || (z >= (-320) + 114880 && z < (-320) + 115200)
							 || (z >= (-320) + 115520 && z < (-320) + 115840)
							 || (z >= (-320) + 116160 && z < (-320) + 116480)
							 || (z >= (-320) + 116800 && z < (-320) + 117120)
							 || (z >= (-320) + 117440 && z < (-320) + 117760)
							 || (z >= (-320) + 118080 && z < (-320) + 118400)
							 || (z >= (-320) + 118720 && z < (-320) + 119040)
							 || (z >= (-320) + 119360 && z < (-320) + 119680)
							 || (z >= (-320) + 120000 && z < (-320) + 120320)
							 || (z >= (-320) + 120640 && z < (-320) + 120960)
							 || (z >= (-320) + 121280 && z < (-320) + 121600)
							 || (z >= (-320) + 121920 && z < (-320) + 122240)
							 || (z >= (-320) + 122560 && z < (-320) + 122880)
							 || (z >= (-320) + 123200 && z < (-320) + 123520)
							 || (z >= (-320) + 123840 && z < (-320) + 124160)
							 || (z >= (-320) + 124480 && z < (-320) + 124800)
							 || (z >= (-320) + 125120 && z < (-320) + 125440)
							 || (z >= (-320) + 125760 && z < (-320) + 126080)
							 || (z >= (-320) + 126040 && z < (-320) + 126720)
							 || (z >= (-320) + 127040 && z < (-320) + 127360)
							 || (z >= (-320) + 127680 && z < (-320) + 128000)
							 || (z >= (-320) + 128320 && z < (-320) + 128640)
							 || (z >= (-320) + 128960 && z < (-320) + 129280)
							 || (z >= (-320) + 129600 && z < (-320) + 129920)
							 || (z >= (-320) + 130240 && z < (-320) + 130560)
							 || (z >= (-320) + 130880 && z < (-320) + 131200)
							 || (z >= (-320) + 131520 && z < (-320) + 131840)
							 || (z >= (-320) + 132160 && z < (-320) + 132480)
							 || (z >= (-320) + 132800 && z < (-320) + 133120)
							 || (z >= (-320) + 133440 && z < (-320) + 133760)
							 || (z >= (-320) + 134080 && z < (-320) + 134400)
							 || (z >= (-320) + 134720 && z < (-320) + 135040)
							 || (z >= (-320) + 135360 && z < (-320) + 135680)
							 || (z >= (-320) + 136000 && z < (-320) + 136320)
							 || (z >= (-320) + 136640 && z < (-320) + 136960)
							 || (z >= (-320) + 137280 && z < (-320) + 137600)
							 || (z >= (-320) + 137920 && z < (-320) + 138240)
							 || (z >= (-320) + 138560 && z < (-320) + 138880)
							 || (z >= (-320) + 139200 && z < (-320) + 139520)
							 || (z >= (-320) + 139840 && z < (-320) + 140160)
							 || (z >= (-320) + 140480 && z < (-320) + 140800)
							 || (z >= (-320) + 141121 && z < (-320) + 141440)
							 || (z >= (-320) + 141760 && z < (-320) + 142080)
							 || (z >= (-320) + 142400 && z < (-320) + 142720)
							 || (z >= (-320) + 143040 && z < (-320) + 143360)
							 || (z >= (-320) + 143680 && z < (-320) + 144000)
							 || (z >= (-320) + 144320 && z < (-320) + 144640)
							 || (z >= (-320) + 144960 && z < (-320) + 145280)
							 || (z >= (-320) + 145600 && z < (-320) + 145920)
							 || (z >= (-320) + 146240 && z < (-320) + 146560)
							 || (z >= (-320) + 146880 && z < (-320) + 147200)
							 || (z >= (-320) + 147520 && z < (-320) + 147840)
							 || (z >= (-320) + 148160 && z < (-320) + 148480)
							 || (z >= (-320) + 148800 && z < (-320) + 149120)
							 || (z >= (-320) + 149440 && z < (-320) + 149760)
							 || (z >= (-320) + 150080 && z < (-320) + 150400)
							 || (z >= (-320) + 150720 && z < (-320) + 151040)
							 || (z >= (-320) + 151360 && z < (-320) + 151680)
							 || (z >= (-320) + 152000 && z < (-320) + 152320)
							 || (z >= (-320) + 152640 && z < (-320) + 152960)
							 || (z >= (-320) + 153280 && z < (-320) + 153600)
							 || (z >= (-320) + 153920 && z < (-320) + 154240)
							 || (z >= (-320) + 154560 && z < (-320) + 154880)
							 || (z >= (-320) + 155200 && z < (-320) + 155520)
							 || (z >= (-320) + 155840 && z < (-320) + 156160)
							 || (z >= (-320) + 156480 && z < (-320) + 156800)
							 || (z >= (-320) + 157120 && z < (-320) + 157440)
							 || (z >= (-320) + 157760 && z < (-320) + 158080)
							 || (z >= (-320) + 158400 && z < (-320) + 158720)
							 || (z >= (-320) + 159040 && z < (-320) + 159360)
							 || (z >= (-320) + 159680 && z < (-320) + 160000)
							 || (z >= (-320) + 160320 && z < (-320) + 160640)
							 || (z >= (-320) + 160960 && z < (-320) + 161280)
							 || (z >= (-320) + 161600 && z < (-320) + 161920)
							 || (z >= (-320) + 162240 && z < (-320) + 162560)
							 || (z >= (-320) + 162880 && z < (-320) + 163200)
							 || (z >= (-320) + 163520 && z < (-320) + 163840)
							 || (z >= (-320) + 164160 && z < (-320) + 164480)
							 || (z >= (-320) + 164800 && z < (-320) + 165120)
							 || (z >= (-320) + 165440 && z < (-320) + 165760)
							 || (z >= (-320) + 166080 && z < (-320) + 166400)
							 || (z >= (-320) + 166720 && z < (-320) + 167040)
							 || (z >= (-320) + 167360 && z < (-320) + 167680)
							 || (z >= (-320) + 168000 && z < (-320) + 168320)
							 || (z >= (-320) + 168640 && z < (-320) + 168960)
							 || (z >= (-320) + 169280 && z < (-320) + 169600)
							 || (z >= (-320) + 169920 && z < (-320) + 170240)
							 || (z >= (-320) + 170560 && z < (-320) + 170880)
							 || (z >= (-320) + 171200 && z < (-320) + 171520)
							 || (z >= (-320) + 171840 && z < (-320) + 172160)
							 || (z >= (-320) + 172480 && z < (-320) + 172800)
							 || (z >= (-320) + 173120 && z < (-320) + 173440)
							 || (z >= (-320) + 173760 && z < (-320) + 174080)
							 || (z >= (-320) + 174400 && z < (-320) + 174720)
							 || (z >= (-320) + 175040 && z < (-320) + 175360)
							 || (z >= (-320) + 175680 && z < (-320) + 176000)
							 || (z >= (-320) + 176320 && z < (-320) + 176640)
							 || (z >= (-320) + 176960 && z < (-320) + 177280)
							 || (z >= (-320) + 177600 && z < (-320) + 177920)
							 || (z >= (-320) + 178240 && z < (-320) + 178560)
							 || (z >= (-320) + 178880 && z < (-320) + 179200)
							 || (z >= (-320) + 179520 && z < (-320) + 179840)
							 || (z >= (-320) + 180160 && z < (-320) + 180480)
							 || (z >= (-320) + 180800 && z < (-320) + 181120)
							 || (z >= (-320) + 181440 && z < (-320) + 181760)
							 || (z >= (-320) + 182080 && z < (-320) + 182400)
							 || (z >= (-320) + 182720 && z < (-320) + 183040)
							 || (z >= (-320) + 183360 && z < (-320) + 183680)
							 || (z >= (-320) + 184000 && z < (-320) + 184320)
							 || (z >= (-320) + 184640 && z < (-320) + 184960)
							 || (z >= (-320) + 185280 && z < (-320) + 185600)
							 || (z >= (-320) + 185920 && z < (-320) + 186240)
							 || (z >= (-320) + 186560 && z < (-320) + 186880)
							 || (z >= (-320) + 187200 && z < (-320) + 187520)
							 || (z >= (-320) + 187840 && z < (-320) + 188160)
							 || (z >= (-320) + 188480 && z < (-320) + 188800)
							 || (z >= (-320) + 189120 && z < (-320) + 189440)
							 || (z >= (-320) + 189760 && z < (-320) + 190080)
							 || (z >= (-320) + 190400 && z < (-320) + 190720)
							 || (z >= (-320) + 191040 && z < (-320) + 191360)
							 || (z >= (-320) + 191680 && z < (-320) + 192000)
							 || (z >= (-320) + 192320 && z < (-320) + 192640)
							 || (z >= (-320) + 192960 && z < (-320) + 193280)
							 || (z >= (-320) + 193600 && z < (-320) + 193920)
							 || (z >= (-320) + 194240 && z < (-320) + 194560)
							 || (z >= (-320) + 194880 && z < (-320) + 195200)
							 || (z >= (-320) + 195520 && z < (-320) + 195840)
							 || (z >= (-320) + 196160 && z < (-320) + 196480)
							 || (z >= (-320) + 196800 && z < (-320) + 197120)
							 || (z >= (-320) + 197440 && z < (-320) + 197760)
							 || (z >= (-320) + 198080 && z < (-320) + 198400)
							 || (z >= (-320) + 198720 && z < (-320) + 199040)
							 || (z >= (-320) + 199360 && z < (-320) + 199680)
							 || (z >= (-320) + 200000 && z < (-320) + 200320)
							 || (z >= (-320) + 200640 && z < (-320) + 200960)
							 || (z >= (-320) + 201280 && z < (-320) + 201600)
							 || (z >= (-320) + 201920 && z < (-320) + 202240)
							 || (z >= (-320) + 202560 && z < (-320) + 202880)
							 || (z >= (-320) + 203200 && z < (-320) + 203520)
							 || (z >= (-320) + 203840 && z < (-320) + 204160)
							 || (z >= (-320) + 204480 && z < (-320) + 204800)
							 || (z >= (-320) + 205120 && z < (-320) + 205440)
							 || (z >= (-320) + 205760 && z < (-320) + 206080)
							 || (z >= (-320) + 206400 && z < (-320) + 206720)
							 || (z >= (-320) + 207040 && z < (-320) + 207360)
							 || (z >= (-320) + 207680 && z < (-320) + 208000)
							 || (z >= (-320) + 208320 && z < (-320) + 208640)
							 || (z >= (-320) + 208960 && z < (-320) + 209280)
							 || (z >= (-320) + 209600 && z < (-320) + 209320)
							 || (z >= (-320) + 210240 && z < (-320) + 210560)
							 || (z >= (-320) + 210880 && z < (-320) + 211200)
							 || (z >= (-320) + 211520 && z < (-320) + 211840)
							 || (z >= (-320) + 212160 && z < (-320) + 212480)
							 || (z >= (-320) + 212800 && z < (-320) + 213120)
							 || (z >= (-320) + 213440 && z < (-320) + 213760)
							 || (z >= (-320) + 214080 && z < (-320) + 214400)
							 || (z >= (-320) + 214720 && z < (-320) + 215040)
							 || (z >= (-320) + 215360 && z < (-320) + 215680)
							 || (z >= (-320) + 216000 && z < (-320) + 216320)
							 || (z >= (-320) + 216640 && z < (-320) + 216960)
							 || (z >= (-320) + 217280 && z < (-320) + 217600)
							 || (z >= (-320) + 217920 && z < (-320) + 218240)
							 || (z >= (-320) + 218560 && z < (-320) + 218880)
							 || (z >= (-320) + 219200 && z < (-320) + 219520)
							 || (z >= (-320) + 219840 && z < (-320) + 220160)
							 || (z >= (-320) + 220480 && z < (-320) + 220800)
							 || (z >= (-320) + 221120 && z < (-320) + 221440)
							 || (z >= (-320) + 221760 && z < (-320) + 222080)
							 || (z >= (-320) + 222400 && z < (-320) + 222720)
							 || (z >= (-320) + 223040 && z < (-320) + 223360)
							 || (z >= (-320) + 223680 && z < (-320) + 224000)
							 || (z >= (-320) + 224320 && z < (-320) + 224640)
							 || (z >= (-320) + 224960 && z < (-320) + 225280)
							 || (z >= (-320) + 225600 && z < (-320) + 225920)
							 || (z >= (-320) + 226240 && z < (-320) + 226560)
							 || (z >= (-320) + 226880 && z < (-320) + 227200)
							 || (z >= (-320) + 227520 && z < (-320) + 227840)
							 || (z >= (-320) + 228160 && z < (-320) + 228480)
							 || (z >= (-320) + 228800 && z < (-320) + 229120)
							 || (z >= (-320) + 229440 && z < (-320) + 229760)
							 || (z >= (-320) + 230080 && z < (-320) + 230400)
							 || (z >= (-320) + 230720 && z < (-320) + 231040)
							 || (z >= (-320) + 231360 && z < (-320) + 231680)
							 || (z >= (-320) + 232000 && z < (-320) + 232320)
							 || (z >= (-320) + 232640 && z < (-320) + 232960)
							 || (z >= (-320) + 233280 && z < (-320) + 233600)
							 || (z >= (-320) + 233920 && z < (-320) + 234240)
							 || (z >= (-320) + 234560 && z < (-320) + 234880)
							 || (z >= (-320) + 235200 && z < (-320) + 235520)
							 || (z >= (-320) + 235840 && z < (-320) + 236160)
							 || (z >= (-320) + 236480 && z < (-320) + 236800)
							 || (z >= (-320) + 237120 && z < (-320) + 237440)
							 || (z >= (-320) + 237760 && z < (-320) + 238080)
							 || (z >= (-320) + 238400 && z < (-320) + 238720)
							 || (z >= (-320) + 239040 && z < (-320) + 239360)
							 || (z >= (-320) + 239680 && z < (-320) + 240000)
							 || (z >= (-320) + 240320 && z < (-320) + 240640)
							 || (z >= (-320) + 240960 && z < (-320) + 241280)
							 || (z >= (-320) + 241600 && z < (-320) + 241920)
							 || (z >= (-320) + 242240 && z < (-320) + 242560)
							 || (z >= (-320) + 242880 && z < (-320) + 243200)
							 || (z >= (-320) + 243520 && z < (-320) + 243840)
							 || (z >= (-320) + 244160 && z < (-320) + 244480)
							 || (z >= (-320) + 244800 && z < (-320) + 245120)
							 || (z >= (-320) + 245440 && z < (-320) + 245760)
							 || (z >= (-320) + 246080 && z < (-320) + 246400)
							 || (z >= (-320) + 246720 && z < (-320) + 247040)
							 || (z >= (-320) + 247360 && z < (-320) + 247680)
							 || (z >= (-320) + 248000 && z < (-320) + 248320)
							 || (z >= (-320) + 248640 && z < (-320) + 248960)
							 || (z >= (-320) + 249280 && z < (-320) + 249600)
							 || (z >= (-320) + 249920 && z < (-320) + 250240)
							 || (z >= (-320) + 250560 && z < (-320) + 250880)
							 || (z >= (-320) + 251200 && z < (-320) + 251520)
							 || (z >= (-320) + 251840 && z < (-320) + 252160)
							 || (z >= (-320) + 252480 && z < (-320) + 252800)
							 || (z >= (-320) + 253120 && z < (-320) + 253440)
							 || (z >= (-320) + 253760 && z < (-320) + 254080)
							 || (z >= (-320) + 254400 && z < (-320) + 254720)
							 || (z >= (-320) + 255040 && z < (-320) + 255360)
							 || (z >= (-320) + 255680 && z < (-320) + 256000)
							 || (z >= (-320) + 256320 && z < (-320) + 256640)
							 || (z >= (-320) + 256960 && z < (-320) + 257280)
							 || (z >= (-320) + 257600 && z < (-320) + 257920)
							 || (z >= (-320) + 258240 && z < (-320) + 258560)
							 || (z >= (-320) + 258880 && z < (-320) + 259200)
							 || (z >= (-320) + 259520 && z < (-320) + 259840)
							 || (z >= (-320) + 260160 && z < (-320) + 260480)
							 || (z >= (-320) + 260800 && z < (-320) + 261120)
							 || (z >= (-320) + 261440 && z < (-320) + 261760)
							 || (z >= (-320) + 262080 && z < (-320) + 262400)
							 || (z >= (-320) + 262720 && z < (-320) + 263040)
							 || (z >= (-320) + 263360 && z < (-320) + 236680)
							 || (z >= (-320) + 264000 && z < (-320) + 264320)
							 || (z >= (-320) + 264640 && z < (-320) + 264960)
							 || (z >= (-320) + 265280 && z < (-320) + 265600)
							 || (z >= (-320) + 265920 && z < (-320) + 266240)
							 || (z >= (-320) + 266560 && z < (-320) + 266880)
							 || (z >= (-320) + 267200 && z < (-320) + 267520)
							 || (z >= (-320) + 267840 && z < (-320) + 268160)
							 || (z >= (-320) + 268480 && z < (-320) + 268800)
							 || (z >= (-320) + 269120 && z < (-320) + 269440)
							 || (z >= (-320) + 269760 && z < (-320) + 270080)
							 || (z >= (-320) + 270400 && z < (-320) + 270720)
							 || (z >= (-320) + 271040 && z < (-320) + 271360)
							 || (z >= (-320) + 271680 && z < (-320) + 272000)
							 || (z >= (-320) + 272320 && z < (-320) + 272640)
							 || (z >= (-320) + 272960 && z < (-320) + 273280)
							 || (z >= (-320) + 273600 && z < (-320) + 273920)
							 || (z >= (-320) + 272240 && z < (-320) + 274560)
							 || (z >= (-320) + 274880 && z < (-320) + 275200)
							 || (z >= (-320) + 275520 && z < (-320) + 275840)
							 || (z >= (-320) + 276160 && z < (-320) + 276480)
							 || (z >= (-320) + 276800 && z < (-320) + 277120)
							 || (z >= (-320) + 277440 && z < (-320) + 277760)
							 || (z >= (-320) + 278080 && z < (-320) + 278400)
							 || (z >= (-320) + 278720 && z < (-320) + 279040)
							 || (z >= (-320) + 279360 && z < (-320) + 279680)
							 || (z >= (-320) + 280000 && z < (-320) + 280320)
							 || (z >= (-320) + 280640 && z < (-320) + 280960)
							 || (z >= (-320) + 281280 && z < (-320) + 281600)
							 || (z >= (-320) + 281920 && z < (-320) + 282240)
							 || (z >= (-320) + 282560 && z < (-320) + 282880)
							 || (z >= (-320) + 283200 && z < (-320) + 283520)
							 || (z >= (-320) + 283840 && z < (-320) + 284160)
							 || (z >= (-320) + 284480 && z < (-320) + 284800)
							 || (z >= (-320) + 285120 && z < (-320) + 285440)
							 || (z >= (-320) + 285760 && z < (-320) + 286080)
							 || (z >= (-320) + 286400 && z < (-320) + 286720)
							 || (z >= (-320) + 287040 && z < (-320) + 287360)
							 || (z >= (-320) + 287680 && z < (-320) + 288000)
							 || (z >= (-320) + 288320 && z < (-320) + 288640)
							 || (z >= (-320) + 288960 && z < (-320) + 289280)
							 || (z >= (-320) + 289600 && z < (-320) + 289920)
							 || (z >= (-320) + 290240 && z < (-320) + 290560)
							 || (z >= (-320) + 290880 && z < (-320) + 291200)
							 || (z >= (-320) + 291520 && z < (-320) + 291840)
							 || (z >= (-320) + 292160 && z < (-320) + 292480)
							 || (z >= (-320) + 292800 && z < (-320) + 293120)
							 || (z >= (-320) + 293440 && z < (-320) + 293760)
							 || (z >= (-320) + 294080 && z < (-320) + 294400)
							 || (z >= (-320) + 294720 && z < (-320) + 295040)
							 || (z >= (-320) + 295360 && z < (-320) + 295680)
							 || (z >= (-320) + 296000 && z < (-320) + 296320)
							 || (z >= (-320) + 296640 && z < (-320) + 296960)
							 || (z >= (-320) + 297280 && z < (-320) + 297600)
							 || (z >= (-320) + 297920 && z < (-320) + 298240)
							 || (z >= (-320) + 298560 && z < (-320) + 298880)
							 || (z >= (-320) + 299200 && z < (-320) + 299520)
							 || (z >= (-320) + 299840 && z < (-320) + 300160)
							 || (z >= (-320) + 300480 && z < (-320) + 300800)
							 || (z >= (-320) + 301120 && z < (-320) + 301440)
							 || (z >= (-320) + 301760 && z < (-320) + 302080)
							 || (z >= (-320) + 302400 && z < (-320) + 302720)
							 || (z >= (-320) + 303040 && z < (-320) + 303360)
							 || (z >= (-320) + 303680 && z < (-320) + 304000)
							 || (z >= (-320) + 304320 && z < (-320) + 304640)
							 || (z >= (-320) + 304960 && z < (-320) + 305280)
							 || (z >= (-320) + 305600 && z < (-320) + 305920)
							 || (z >= (-320) + 306240 && z < (-320) + 306560)
							 || (z >= (-320) + 306880 && z < (-320) + 307200))
						begin
						//This is executed when the white pixel belongs to the left half(c direction)
							c = c+1;
						end
						if(z >= 152960 && z < 307200)
						begin
						//This is executed when the white pixel belongs to the bottom half(d direction)
							d=d+1;
						end
					end
					z = z + 1;
					//We increment z after looking at every pixel so that we can keep track of the pixels we have read
			end
			if(k==0)
			begin
			//We execute the algorithm when k = 0(ie. when we have finished reading a frame
			end
		end
		algorithmtester U1 (a, b, c, d, k, LEDR);
endmodule